module AND2(
    input  wire A,
    input  wire B,
    output wire Y
);

   and _and2(Y, A, B);

endmodule
