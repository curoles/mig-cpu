module TbTop (
    input  wire clk
    //input  wire [WIDTH-1:0]  in,
    //input  wire              en,
    //output wire [SIZE-1:0]   out
);


    ///*output  reg*/ wire [6:0]  opcode;
    ///*output  reg*/ wire [4:0]  rd, rs1, rs2;
    ///*output  reg*/ wire [2:0]  funct3;
    ///*output  reg*/ wire [6:0]  funct7;
    ///*output  reg*/ wire [31:0] imm;

    //RiscvInsnTypeDecode _insn_type_decode(
    //    .clk(clk), .insn(insn),
    //    .opcode(opcode),
    //    .rd(rd), .rs1(rs1), .rs2(rs2),
    //    .funct3(funct3), .funct7(funct7),
    //    .imm(imm)
    //);

endmodule : TbTop
