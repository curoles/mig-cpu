/* 3-inputs NAND gate.
 *
 *
 * http://bibl.ica.jku.at/dc/build/html/basiccircuits/basiccircuits.html
 */
